-- #P7i6 ULA 
-- EDUARDO A. MARRAS DE SOUZA RA: 20078408
-- BIANCA A. ANDRADE RA: 21007245
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY ULA IS
PORT ( A, B : IN  STD_LOGIC_VECTOR(7 DOWNTO 0) ; -- DUAS ENTRADAS PARA OPERAÇÃO
ADDSUBC : IN STD_LOGIC; -- CONTROLADOR DE OPERAÇÃO (ADD OU SUB)
S  : OUT  STD_LOGIC_VECTOR(7 DOWNTO 0) ) ; -- SAÍDA DA ULA
END ULA ;

ARCHITECTURE LOGIC OF ULA IS    
BEGIN
S <= A + B WHEN ADDSUBC = '0' ELSE A + (NOT B) + 1; -- QUANDO CONTROLADOR FOR 0, SOMA. QUANDO FOR 1, SUBTRAÇÃO.
END LOGIC ;