-- #P7i6 REGISTRADOR
-- EDUARDO A. MARRAS DE SOUZA RA: 20078408
-- BIANCA A. ANDRADE RA: 21007245
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY REG IS
PORT (  D : IN  STD_LOGIC_VECTOR(7 DOWNTO 0) ; -- ENTRADA DO REGISTRADOR
RIN, CLOCK : IN  STD_LOGIC ; -- ENTRADA PARA O ENABLE E ENTRADA PARA O CLOCK DO REGISTRADOR
Q  : OUT  STD_LOGIC_VECTOR(7 DOWNTO 0) ) ; -- SAÍDA DO REGISTRADOR
END REG ;

ARCHITECTURE LOGIC OF REG IS
BEGIN
PROCESS ( CLOCK ) -- PROCESSO EM FUNÇÃO DO CLOCK
BEGIN
IF RIN = '1' THEN -- SE O ENABLE FOR ATIVADO
IF CLOCK'EVENT AND CLOCK = '1' THEN -- SE O CLOCK SUBIR
Q <= D ; -- SAÍDA RECEBE A ENTRADA
END IF ;
END IF;
END PROCESS ;
END LOGIC ;