-- #P7i6 - DATA H
-- EDUARDO A. MARRAS DE SOUZA RA: 20078408
-- BIANCA A. ANDRADE RA: 21007245
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY DATA IS

PORT (CLOCK, R0IN, R0T, R1IN, R1T, R2IN, R2T, R3IN, R3T, AIN, GIN, GOUT, ADDSUB, EXTERN : IN STD_LOGIC; -- ENTRADAS SIMPLES DO DATA
		DATAENT : IN STD_LOGIC_VECTOR(7 DOWNTO 0); -- ENTRADA DE DATA DO CIRCUITO, COM 8 BITS
		BARRAMENTO : INOUT STD_LOGIC_VECTOR(7 DOWNTO 0) ); -- BARRAMENTO DO TIPO INOUT COM 8 BITS PARA ENVIO E RECEBIMENTO DE DADOS
END DATA;


ARCHITECTURE LOGIC OF DATA IS    
SIGNAL AS, RES, GS, R0S, R1S, R2S, R3S: STD_LOGIC_VECTOR(7 DOWNTO 0); -- SINAIS PARA O DATA

COMPONENT REG -- DECLARAÇÃO DOS COMPONENTES

PORT(D : IN  STD_LOGIC_VECTOR(7 DOWNTO 0);
RIN, CLOCK : IN  STD_LOGIC ;
Q  : OUT  STD_LOGIC_VECTOR(7 DOWNTO 0));

END COMPONENT ;

COMPONENT ULA 

PORT (A, B : IN  STD_LOGIC_VECTOR(7 DOWNTO 0) ;
ADDSUBC : IN STD_LOGIC;
S  : OUT  STD_LOGIC_VECTOR(7 DOWNTO 0) ) ;

END COMPONENT;

COMPONENT TRISTATE 
PORT (INPUT : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
            ENABLE: IN STD_LOGIC;
            OUTPUT     : OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END COMPONENT;

BEGIN -- PORT MAPS DOS COMPONENTES LISTADOS

R0: REG PORT MAP(BARRAMENTO, R0IN, CLOCK, R0S);
R1: REG PORT MAP(BARRAMENTO, R1IN, CLOCK, R1S);
R2: REG PORT MAP(BARRAMENTO, R2IN, CLOCK, R2S);
R3: REG PORT MAP(BARRAMENTO, R3IN, CLOCK, R3S);
A: REG PORT MAP(BARRAMENTO, AIN, CLOCK, AS);
G: REG PORT MAP(RES, GIN, CLOCK, GS);

TRG: TRISTATE PORT MAP(GS, GOUT, BARRAMENTO);
TRD: TRISTATE PORT MAP(DATAENT, EXTERN, BARRAMENTO);
TR0: TRISTATE PORT MAP(R0S, R0T, BARRAMENTO);
TR1: TRISTATE PORT MAP(R1S, R1T, BARRAMENTO);
TR2: TRISTATE PORT MAP(R2S, R2T, BARRAMENTO);
TR3: TRISTATE PORT MAP(R3S, R3T, BARRAMENTO);

UL: ULA PORT MAP(AS, BARRAMENTO, ADDSUB, RES);

END LOGIC ;